magic
tech sky130A
timestamp 1736697198
<< nwell >>
rect -905 -13 -595 149
rect -115 -12 224 133
rect -903 -14 -617 -13
<< nmos >>
rect -351 -160 -336 -115
rect -48 -164 -33 -122
rect 108 -160 123 -118
rect -794 -299 -779 -257
rect -69 -411 -54 -368
<< pmos >>
rect -794 26 -779 68
rect -48 9 -33 51
rect 108 11 123 56
<< ndiff >>
rect -398 -128 -351 -115
rect -398 -147 -379 -128
rect -362 -147 -351 -128
rect -398 -160 -351 -147
rect -336 -128 -289 -115
rect -336 -147 -320 -128
rect -303 -147 -289 -128
rect -336 -160 -289 -147
rect -92 -134 -48 -122
rect -92 -152 -81 -134
rect -64 -152 -48 -134
rect -92 -164 -48 -152
rect -33 -132 8 -122
rect -33 -150 -19 -132
rect -2 -150 8 -132
rect -33 -164 8 -150
rect 74 -131 108 -118
rect 74 -149 81 -131
rect 98 -149 108 -131
rect 74 -160 108 -149
rect 123 -129 176 -118
rect 123 -147 136 -129
rect 153 -147 176 -129
rect 123 -160 176 -147
rect -831 -270 -794 -257
rect -831 -287 -826 -270
rect -809 -287 -794 -270
rect -831 -299 -794 -287
rect -779 -269 -727 -257
rect -779 -286 -756 -269
rect -739 -286 -727 -269
rect -779 -299 -727 -286
rect -106 -379 -69 -368
rect -106 -398 -94 -379
rect -76 -398 -69 -379
rect -106 -411 -69 -398
rect -54 -379 1 -368
rect -54 -398 -38 -379
rect -20 -398 1 -379
rect -54 -411 1 -398
<< pdiff >>
rect -828 56 -794 68
rect -828 39 -821 56
rect -804 39 -794 56
rect -828 26 -794 39
rect -779 57 -724 68
rect -779 40 -756 57
rect -739 40 -724 57
rect -779 26 -724 40
rect -90 40 -48 51
rect -90 22 -82 40
rect -65 22 -48 40
rect -90 9 -48 22
rect -33 41 10 51
rect -33 23 -15 41
rect 2 23 10 41
rect -33 9 10 23
rect 68 43 108 56
rect 68 25 79 43
rect 96 25 108 43
rect 68 11 108 25
rect 123 42 170 56
rect 123 24 143 42
rect 160 24 170 42
rect 123 11 170 24
<< ndiffc >>
rect -379 -147 -362 -128
rect -320 -147 -303 -128
rect -81 -152 -64 -134
rect -19 -150 -2 -132
rect 81 -149 98 -131
rect 136 -147 153 -129
rect -826 -287 -809 -270
rect -756 -286 -739 -269
rect -94 -398 -76 -379
rect -38 -398 -20 -379
<< pdiffc >>
rect -821 39 -804 56
rect -756 40 -739 57
rect -82 22 -65 40
rect -15 23 2 41
rect 79 25 96 43
rect 143 24 160 42
<< psubdiff >>
rect 48 -194 184 -193
rect -90 -196 184 -194
rect -90 -213 -38 -196
rect -17 -199 184 -196
rect -17 -213 13 -199
rect -90 -216 13 -213
rect 34 -216 123 -199
rect 144 -216 184 -199
rect -90 -218 184 -216
rect -415 -235 -284 -231
rect -415 -237 -332 -235
rect -415 -254 -403 -237
rect -382 -252 -332 -237
rect -311 -252 -284 -235
rect -382 -254 -284 -252
rect -415 -258 -284 -254
rect -836 -354 -705 -344
rect -836 -384 -778 -354
rect -756 -355 -705 -354
rect -756 -384 -739 -355
rect -836 -385 -739 -384
rect -717 -385 -705 -355
rect -836 -395 -705 -385
rect -112 -485 -12 -483
rect -112 -486 -49 -485
rect -112 -503 -99 -486
rect -79 -502 -49 -486
rect -29 -502 -12 -485
rect -79 -503 -12 -502
rect -112 -507 -12 -503
<< nsubdiff >>
rect -886 122 -624 124
rect -886 120 -670 122
rect -886 101 -745 120
rect -719 103 -670 120
rect -644 103 -624 122
rect -719 101 -624 103
rect -886 97 -624 101
rect -94 108 167 110
rect -94 91 -34 108
rect -15 91 13 108
rect 32 107 167 108
rect 32 91 114 107
rect -94 90 114 91
rect 133 90 167 107
rect -94 86 167 90
<< psubdiffcont >>
rect -38 -213 -17 -196
rect 13 -216 34 -199
rect 123 -216 144 -199
rect -403 -254 -382 -237
rect -332 -252 -311 -235
rect -778 -384 -756 -354
rect -739 -385 -717 -355
rect -99 -503 -79 -486
rect -49 -502 -29 -485
<< nsubdiffcont >>
rect -745 101 -719 120
rect -670 103 -644 122
rect -34 91 -15 108
rect 13 91 32 108
rect 114 90 133 107
<< poly >>
rect -794 68 -779 85
rect -48 51 -33 64
rect 108 56 123 70
rect -794 -58 -779 26
rect -48 -42 -33 9
rect -862 -59 -779 -58
rect -874 -79 -779 -59
rect -92 -47 -33 -42
rect 108 -47 123 11
rect -92 -64 -84 -47
rect -62 -64 -33 -47
rect -92 -70 -33 -64
rect -874 -96 -837 -79
rect -817 -96 -779 -79
rect -874 -109 -779 -96
rect -865 -110 -779 -109
rect -794 -257 -779 -110
rect -351 -115 -336 -101
rect -48 -122 -33 -70
rect 68 -56 123 -47
rect 68 -73 85 -56
rect 107 -73 123 -56
rect 68 -80 123 -73
rect 79 -81 123 -80
rect 108 -118 123 -81
rect -351 -176 -336 -160
rect -387 -181 -336 -176
rect -387 -198 -379 -181
rect -359 -198 -336 -181
rect -48 -188 -33 -164
rect 108 -182 123 -160
rect -387 -203 -336 -198
rect -351 -224 -336 -203
rect -794 -329 -779 -299
rect -69 -368 -54 -336
rect -69 -424 -54 -411
rect -109 -432 -54 -424
rect -109 -449 -97 -432
rect -77 -449 -54 -432
rect -109 -455 -54 -449
rect -69 -463 -54 -455
<< polycont >>
rect -84 -64 -62 -47
rect -837 -96 -817 -79
rect 85 -73 107 -56
rect -379 -198 -359 -181
rect -97 -449 -77 -432
<< locali >>
rect -979 213 -932 214
rect -560 213 -528 215
rect -979 189 -527 213
rect -979 -55 -932 189
rect -561 170 -528 189
rect -561 145 -529 170
rect -886 122 -624 124
rect -886 120 -670 122
rect -886 101 -823 120
rect -797 101 -745 120
rect -719 103 -670 120
rect -644 103 -624 122
rect -719 101 -624 103
rect -886 97 -624 101
rect -826 64 -796 97
rect -827 56 -795 64
rect -827 39 -821 56
rect -804 39 -795 56
rect -827 30 -795 39
rect -763 57 -731 65
rect -763 40 -756 57
rect -739 40 -731 57
rect -763 31 -731 40
rect -979 -79 -789 -55
rect -979 -96 -837 -79
rect -817 -96 -789 -79
rect -979 -107 -789 -96
rect -946 -110 -789 -107
rect -762 -90 -731 31
rect -762 -92 -616 -90
rect -762 -121 -615 -92
rect -762 -158 -728 -121
rect -649 -158 -615 -121
rect -831 -270 -800 -256
rect -831 -287 -826 -270
rect -809 -287 -800 -270
rect -831 -298 -800 -287
rect -832 -344 -800 -298
rect -762 -269 -731 -158
rect -762 -286 -756 -269
rect -739 -286 -731 -269
rect -762 -299 -731 -286
rect -836 -354 -705 -344
rect -836 -355 -778 -354
rect -836 -385 -826 -355
rect -804 -384 -778 -355
rect -756 -355 -705 -354
rect -756 -384 -739 -355
rect -804 -385 -739 -384
rect -717 -385 -705 -355
rect -836 -395 -705 -385
rect -645 -424 -615 -158
rect -560 -181 -530 145
rect -94 108 167 110
rect -94 107 -34 108
rect -94 90 -84 107
rect -65 91 -34 107
rect -15 91 13 108
rect 32 107 167 108
rect 32 91 78 107
rect -65 90 78 91
rect 97 90 114 107
rect 133 90 167 107
rect -94 86 167 90
rect -89 40 -57 86
rect 74 56 104 86
rect -89 22 -82 40
rect -65 22 -57 40
rect -89 13 -57 22
rect -23 41 9 49
rect -23 23 -15 41
rect 2 23 9 41
rect -330 -47 -48 -41
rect -330 -64 -84 -47
rect -62 -64 -48 -47
rect -387 -128 -353 -67
rect -330 -70 -48 -64
rect -23 -46 9 23
rect 73 43 104 56
rect 73 25 79 43
rect 96 25 104 43
rect 73 14 104 25
rect 137 42 167 55
rect 137 24 143 42
rect 160 24 167 42
rect 137 14 167 24
rect 137 -45 166 14
rect 226 -45 304 -44
rect -23 -47 68 -46
rect -23 -56 112 -47
rect -387 -147 -379 -128
rect -362 -147 -353 -128
rect -387 -155 -353 -147
rect -329 -128 -292 -70
rect -329 -147 -320 -128
rect -303 -147 -292 -128
rect -329 -157 -292 -147
rect -389 -177 -351 -176
rect -418 -178 -351 -177
rect -427 -179 -351 -178
rect -496 -181 -351 -179
rect -560 -198 -379 -181
rect -359 -198 -351 -181
rect -560 -203 -351 -198
rect -415 -235 -284 -231
rect -415 -237 -332 -235
rect -415 -254 -403 -237
rect -382 -252 -332 -237
rect -311 -252 -284 -235
rect -382 -254 -284 -252
rect -415 -258 -284 -254
rect -186 -284 -157 -70
rect -23 -73 85 -56
rect 107 -73 112 -56
rect -23 -80 112 -73
rect -23 -124 9 -80
rect 79 -81 111 -80
rect 137 -82 304 -45
rect 137 -83 259 -82
rect 137 -121 166 -83
rect -89 -134 -57 -126
rect -89 -152 -81 -134
rect -64 -152 -57 -134
rect -89 -194 -57 -152
rect -26 -132 6 -124
rect -26 -150 -19 -132
rect -2 -150 6 -132
rect -26 -158 6 -150
rect 78 -131 102 -123
rect 78 -149 81 -131
rect 98 -149 102 -131
rect 78 -159 102 -149
rect 128 -129 166 -121
rect 128 -147 136 -129
rect 153 -147 166 -129
rect 128 -154 166 -147
rect 77 -193 102 -159
rect 48 -194 184 -193
rect -90 -196 184 -194
rect -90 -198 -38 -196
rect -90 -215 -84 -198
rect -63 -213 -38 -198
rect -17 -197 184 -196
rect -17 -199 78 -197
rect -17 -213 13 -199
rect -63 -215 13 -213
rect -90 -216 13 -215
rect 34 -214 78 -199
rect 99 -199 184 -197
rect 99 -214 123 -199
rect 34 -216 123 -214
rect 144 -216 184 -199
rect -90 -218 184 -216
rect 224 -277 259 -83
rect 128 -279 259 -277
rect 81 -280 259 -279
rect -186 -285 -113 -284
rect -186 -306 -70 -285
rect -100 -330 -70 -306
rect -101 -371 -70 -330
rect -47 -299 259 -280
rect -47 -301 229 -299
rect -47 -302 101 -301
rect -102 -379 -71 -371
rect -102 -398 -94 -379
rect -76 -398 -71 -379
rect -102 -407 -71 -398
rect -47 -374 -9 -302
rect -47 -379 -12 -374
rect -47 -398 -38 -379
rect -20 -398 -12 -379
rect -47 -405 -12 -398
rect -47 -406 -15 -405
rect -645 -432 -69 -424
rect -645 -449 -97 -432
rect -77 -449 -69 -432
rect -645 -454 -69 -449
rect -621 -455 -69 -454
rect -621 -457 -140 -455
rect -112 -485 -12 -483
rect -112 -486 -49 -485
rect -112 -503 -99 -486
rect -79 -502 -49 -486
rect -29 -502 -12 -485
rect -79 -503 -12 -502
rect -112 -507 -12 -503
<< viali >>
rect -823 101 -797 120
rect -826 -385 -804 -355
rect -84 90 -65 107
rect 78 90 97 107
rect -84 -215 -63 -198
rect 78 -214 99 -197
<< metal1 >>
rect -886 120 -624 124
rect -886 101 -823 120
rect -797 101 -624 120
rect -886 97 -624 101
rect -94 107 167 110
rect -94 90 -84 107
rect -65 90 78 107
rect 97 90 167 107
rect -94 86 167 90
rect 48 -194 184 -193
rect -90 -197 184 -194
rect -90 -198 78 -197
rect -90 -215 -84 -198
rect -63 -214 78 -198
rect 99 -214 184 -197
rect -63 -215 184 -214
rect -90 -218 184 -215
rect -415 -258 -284 -231
rect -836 -355 -705 -344
rect -836 -385 -826 -355
rect -804 -385 -705 -355
rect -836 -395 -705 -385
rect -112 -507 -12 -483
<< labels >>
flabel locali -372 -86 -372 -86 0 FreeSans 160 0 0 0 D
flabel locali -129 -441 -129 -441 0 FreeSans 80 0 0 0 ~clk
flabel locali 246 -61 246 -61 0 FreeSans 160 0 0 0 OUT
flabel metal1 54 97 54 97 0 FreeSans 80 0 0 0 vdd
flabel metal1 54 -206 54 -206 0 FreeSans 80 0 0 0 gnd
flabel locali -949 -84 -949 -84 0 FreeSans 160 0 0 0 clk
flabel metal1 -858 109 -858 109 0 FreeSans 160 0 0 0 vdd
flabel metal1 -795 -379 -795 -379 0 FreeSans 80 0 0 0 gnd
<< end >>
