magic
tech sky130A
timestamp 1736572094
<< nwell >>
rect -330 328 395 389
rect -332 -63 396 328
<< nmos >>
rect -37 -554 14 -502
<< pmos >>
rect -37 32 14 84
<< ndiff >>
rect -148 -509 -37 -502
rect -148 -550 -113 -509
rect -82 -550 -37 -509
rect -148 -554 -37 -550
rect 14 -509 172 -502
rect 14 -550 105 -509
rect 136 -550 172 -509
rect 14 -554 172 -550
<< pdiff >>
rect -143 76 -37 84
rect -143 45 -127 76
rect -103 45 -37 76
rect -143 32 -37 45
rect 14 77 176 84
rect 14 46 108 77
rect 132 46 176 77
rect 14 32 176 46
<< ndiffc >>
rect -113 -550 -82 -509
rect 105 -550 136 -509
<< pdiffc >>
rect -127 45 -103 76
rect 108 46 132 77
<< psubdiff >>
rect -284 -651 288 -638
rect -284 -733 -271 -651
rect -188 -653 288 -651
rect -188 -733 161 -653
rect -284 -735 161 -733
rect 244 -735 288 -653
rect -284 -742 288 -735
<< nsubdiff >>
rect -254 282 316 297
rect -254 200 -248 282
rect -165 279 316 282
rect -165 200 212 279
rect -254 197 212 200
rect 295 197 316 279
rect -254 179 316 197
<< psubdiffcont >>
rect -271 -733 -188 -651
rect 161 -735 244 -653
<< nsubdiffcont >>
rect -248 200 -165 282
rect 212 197 295 279
<< poly >>
rect -37 84 14 104
rect -37 -199 14 32
rect -117 -210 14 -199
rect -117 -276 -107 -210
rect -51 -276 14 -210
rect -117 -281 14 -276
rect -37 -502 14 -281
rect -37 -604 14 -554
<< polycont >>
rect -107 -276 -51 -210
<< locali >>
rect -254 286 316 297
rect -254 282 -156 286
rect -254 200 -248 282
rect -165 204 -156 282
rect -73 279 316 286
rect -73 204 212 279
rect -165 200 212 204
rect -254 197 212 200
rect 295 197 316 279
rect -254 179 316 197
rect -137 102 -91 179
rect -137 96 -92 102
rect -136 76 -92 96
rect -136 45 -127 76
rect -103 45 -92 76
rect -136 32 -92 45
rect -135 30 -92 32
rect 97 83 143 84
rect 97 77 144 83
rect 97 46 108 77
rect 132 46 144 77
rect -229 -210 -44 -196
rect -229 -276 -107 -210
rect -51 -276 -44 -210
rect -229 -293 -44 -276
rect 97 -199 144 46
rect 97 -281 199 -199
rect -121 -509 -74 -503
rect -121 -550 -113 -509
rect -82 -550 -74 -509
rect -121 -638 -74 -550
rect 97 -509 144 -281
rect 97 -550 105 -509
rect 136 -550 144 -509
rect 97 -554 144 -550
rect -285 -651 290 -638
rect -285 -733 -271 -651
rect -188 -652 290 -651
rect -188 -733 -146 -652
rect -285 -734 -146 -733
rect -63 -653 290 -652
rect -63 -734 161 -653
rect -285 -735 161 -734
rect 244 -735 290 -653
rect -285 -743 290 -735
<< viali >>
rect -156 204 -73 286
rect -146 -734 -63 -652
<< metal1 >>
rect -252 286 318 298
rect -252 204 -156 286
rect -73 204 318 286
rect -252 178 318 204
rect -280 -652 288 -645
rect -280 -734 -146 -652
rect -63 -734 288 -652
rect -280 -738 288 -734
<< labels >>
flabel metal1 22 230 22 230 0 FreeSans 400 0 0 0 vdd
flabel locali -186 -245 -186 -245 0 FreeSans 400 0 0 0 IN
flabel locali 158 -240 158 -240 0 FreeSans 320 0 0 0 OUT
flabel metal1 30 -688 30 -688 0 FreeSans 320 0 0 0 GND
<< end >>
