magic
tech sky130A
timestamp 1736579761
<< nwell >>
rect -98 -22 222 154
<< nmos >>
rect -28 -257 -1 -195
rect 127 -257 153 -195
<< pmos >>
rect -28 -1 -1 57
rect 127 -1 153 57
<< ndiff >>
rect -77 -209 -28 -195
rect -77 -235 -64 -209
rect -46 -235 -28 -209
rect -77 -257 -28 -235
rect -1 -206 127 -195
rect -1 -240 58 -206
rect 82 -240 127 -206
rect -1 -257 127 -240
rect 153 -212 200 -195
rect 153 -238 169 -212
rect 187 -238 200 -212
rect 153 -257 200 -238
<< pdiff >>
rect -76 43 -28 57
rect -76 15 -62 43
rect -45 15 -28 43
rect -76 -1 -28 15
rect -1 -1 127 57
rect 153 44 197 57
rect 153 14 168 44
rect 185 14 197 44
rect 153 -1 197 14
<< ndiffc >>
rect -64 -235 -46 -209
rect 58 -240 82 -206
rect 169 -238 187 -212
<< pdiffc >>
rect -62 15 -45 43
rect 168 14 185 44
<< psubdiff >>
rect -96 -322 223 -309
rect -96 -354 -3 -322
rect 31 -323 223 -322
rect 31 -354 95 -323
rect -96 -355 95 -354
rect 129 -355 223 -323
<< nsubdiff >>
rect -77 129 198 132
rect -77 102 28 129
rect 59 102 126 129
rect 157 102 198 129
rect -77 101 198 102
<< psubdiffcont >>
rect -3 -354 31 -322
rect 95 -355 129 -323
<< nsubdiffcont >>
rect 28 102 59 129
rect 126 102 157 129
<< poly >>
rect -28 57 -1 71
rect 127 57 153 72
rect -28 -77 -1 -1
rect 127 -41 153 -1
rect 91 -47 153 -41
rect 91 -66 100 -47
rect 119 -66 153 -47
rect 91 -71 153 -66
rect -81 -83 -1 -77
rect -81 -102 -66 -83
rect -47 -102 -1 -83
rect -81 -108 -1 -102
rect -28 -195 -1 -108
rect 127 -195 153 -71
rect -28 -295 -1 -257
rect 127 -295 153 -257
<< polycont >>
rect 100 -66 119 -47
rect -66 -102 -47 -83
<< locali >>
rect -81 129 207 132
rect -81 127 28 129
rect -81 104 -65 127
rect -42 104 28 127
rect -81 102 28 104
rect 59 102 126 129
rect 157 102 207 129
rect -81 98 207 102
rect -70 43 -37 98
rect -70 15 -62 43
rect -45 15 -37 43
rect -70 8 -37 15
rect 160 44 193 51
rect 160 14 168 44
rect 185 14 193 44
rect 66 -47 127 -41
rect 66 -66 100 -47
rect 119 -66 127 -47
rect 66 -71 127 -66
rect -124 -83 -29 -75
rect -124 -102 -66 -83
rect -47 -102 -29 -83
rect -124 -108 -29 -102
rect 49 -108 91 -100
rect 49 -137 52 -108
rect 85 -137 91 -108
rect -71 -209 -37 -200
rect -71 -235 -64 -209
rect -46 -235 -37 -209
rect -71 -312 -37 -235
rect 49 -206 91 -137
rect 160 -108 193 14
rect 160 -137 165 -108
rect 188 -137 193 -108
rect 160 -143 193 -137
rect 49 -240 58 -206
rect 82 -240 91 -206
rect 49 -248 91 -240
rect 160 -212 194 -202
rect 160 -238 169 -212
rect 187 -238 194 -212
rect 160 -312 194 -238
rect -92 -322 225 -312
rect -92 -323 -3 -322
rect -92 -352 -68 -323
rect -40 -352 -3 -323
rect -92 -354 -3 -352
rect 31 -323 225 -322
rect 31 -354 95 -323
rect -92 -355 95 -354
rect 129 -352 163 -323
rect 191 -352 225 -323
rect 129 -355 225 -352
rect -92 -358 225 -355
<< viali >>
rect -65 104 -42 127
rect 52 -137 85 -108
rect 165 -137 188 -108
rect -68 -352 -40 -323
rect 163 -352 191 -323
<< metal1 >>
rect -81 127 207 133
rect -81 104 -65 127
rect -42 104 207 127
rect -81 95 207 104
rect 46 -108 271 -100
rect 46 -137 52 -108
rect 85 -137 165 -108
rect 188 -137 271 -108
rect 46 -143 271 -137
rect -87 -323 219 -317
rect -87 -352 -68 -323
rect -40 -352 163 -323
rect 191 -352 219 -323
rect -87 -357 219 -352
<< labels >>
flabel locali -107 -93 -107 -93 0 FreeSans 160 0 0 0 A
flabel locali 73 -59 74 -58 0 FreeSans 160 0 0 0 B
flabel metal1 240 -118 240 -118 0 FreeSans 160 0 0 0 OUT
flabel metal1 60 -338 60 -338 0 FreeSans 80 0 0 0 gnd
flabel metal1 -18 115 -18 115 0 FreeSans 80 0 0 0 vdd
<< end >>
