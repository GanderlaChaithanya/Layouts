magic
tech sky130A
timestamp 1737455450
<< nwell >>
rect -256 129 564 216
rect -255 42 564 129
<< nmos >>
rect -200 -69 -179 -21
rect -62 -106 -42 -60
rect 29 -106 49 -60
rect 210 -109 232 -63
rect 293 -109 315 -63
rect 469 -107 490 -61
<< pmos >>
rect -200 60 -179 108
rect -62 60 -42 104
rect 29 60 49 104
rect 210 64 232 108
rect 293 64 315 108
rect 469 64 490 108
<< ndiff >>
rect -237 -30 -200 -21
rect -237 -58 -231 -30
rect -211 -58 -200 -30
rect -237 -69 -200 -58
rect -179 -30 -143 -21
rect -179 -58 -172 -30
rect -152 -58 -143 -30
rect -179 -69 -143 -58
rect -99 -69 -62 -60
rect -99 -97 -92 -69
rect -72 -97 -62 -69
rect -99 -106 -62 -97
rect -42 -106 29 -60
rect 49 -73 99 -60
rect 49 -101 63 -73
rect 83 -101 99 -73
rect 49 -106 99 -101
rect 167 -72 210 -63
rect 167 -100 175 -72
rect 195 -100 210 -72
rect 167 -109 210 -100
rect 232 -109 293 -63
rect 315 -78 365 -63
rect 315 -97 327 -78
rect 344 -97 365 -78
rect 315 -109 365 -97
rect 421 -70 469 -61
rect 421 -89 431 -70
rect 448 -89 469 -70
rect 421 -107 469 -89
rect 490 -75 533 -61
rect 490 -94 504 -75
rect 521 -94 533 -75
rect 490 -107 533 -94
<< pdiff >>
rect -236 98 -200 108
rect -236 70 -229 98
rect -209 70 -200 98
rect -236 60 -200 70
rect -179 100 -143 108
rect -179 72 -172 100
rect -152 72 -143 100
rect -179 60 -143 72
rect -105 97 -62 104
rect -105 69 -92 97
rect -72 69 -62 97
rect -105 60 -62 69
rect -42 98 29 104
rect -42 70 -22 98
rect -2 70 29 98
rect -42 60 29 70
rect 49 95 95 104
rect 49 67 60 95
rect 80 67 95 95
rect 49 60 95 67
rect 153 97 210 108
rect 153 78 181 97
rect 198 78 210 97
rect 153 64 210 78
rect 232 100 293 108
rect 232 72 253 100
rect 273 72 293 100
rect 232 64 293 72
rect 315 94 366 108
rect 315 75 332 94
rect 349 75 366 94
rect 315 64 366 75
rect 425 96 469 108
rect 425 77 435 96
rect 452 77 469 96
rect 425 64 469 77
rect 490 96 536 108
rect 490 77 506 96
rect 523 77 536 96
rect 490 64 536 77
<< ndiffc >>
rect -231 -58 -211 -30
rect -172 -58 -152 -30
rect -92 -97 -72 -69
rect 63 -101 83 -73
rect 175 -100 195 -72
rect 327 -97 344 -78
rect 431 -89 448 -70
rect 504 -94 521 -75
<< pdiffc >>
rect -229 70 -209 98
rect -172 72 -152 100
rect -92 69 -72 97
rect -22 70 -2 98
rect 60 67 80 95
rect 181 78 198 97
rect 253 72 273 100
rect 332 75 349 94
rect 435 77 452 96
rect 506 77 523 96
<< psubdiff >>
rect 252 -145 552 -143
rect -241 -149 552 -145
rect -241 -150 508 -149
rect -241 -153 240 -150
rect -241 -172 -180 -153
rect -163 -154 -14 -153
rect -163 -172 -102 -154
rect -241 -173 -102 -172
rect -85 -172 -14 -154
rect 3 -169 240 -153
rect 257 -152 508 -150
rect 257 -154 385 -152
rect 257 -169 327 -154
rect 3 -172 327 -169
rect -85 -173 327 -172
rect 344 -171 385 -154
rect 402 -168 508 -152
rect 525 -168 552 -149
rect 402 -171 552 -168
rect 344 -173 552 -171
rect -241 -177 552 -173
rect 252 -178 552 -177
<< nsubdiff >>
rect 248 176 544 177
rect -118 175 544 176
rect -224 174 544 175
rect -224 173 189 174
rect -224 154 -179 173
rect -162 154 -145 173
rect -128 154 -36 173
rect -19 155 189 173
rect 206 155 289 174
rect 306 155 376 174
rect 393 155 495 174
rect 512 155 544 174
rect -19 154 544 155
rect -224 149 544 154
rect -224 148 -116 149
rect 248 148 544 149
<< psubdiffcont >>
rect -180 -172 -163 -153
rect -102 -173 -85 -154
rect -14 -172 3 -153
rect 240 -169 257 -150
rect 327 -173 344 -154
rect 385 -171 402 -152
rect 508 -168 525 -149
<< nsubdiffcont >>
rect -179 154 -162 173
rect -145 154 -128 173
rect -36 154 -19 173
rect 189 155 206 174
rect 289 155 306 174
rect 376 155 393 174
rect 495 155 512 174
<< poly >>
rect -200 108 -179 121
rect -62 104 -42 122
rect 29 104 49 124
rect 210 108 232 126
rect 293 108 315 127
rect 469 108 490 121
rect -200 30 -179 60
rect -62 31 -42 60
rect 29 34 49 60
rect -236 24 -179 30
rect -236 7 -226 24
rect -209 7 -179 24
rect -236 0 -179 7
rect -99 24 -42 31
rect -99 7 -90 24
rect -73 7 -42 24
rect -99 2 -42 7
rect -12 29 49 34
rect 210 30 232 64
rect -12 12 0 29
rect 18 12 49 29
rect -12 3 49 12
rect -200 -21 -179 0
rect -62 -60 -42 2
rect 29 -60 49 3
rect 169 23 232 30
rect 169 6 185 23
rect 203 6 232 23
rect 169 0 232 6
rect -200 -100 -179 -69
rect 210 -63 232 0
rect 293 33 315 64
rect 293 26 356 33
rect 293 9 321 26
rect 339 9 356 26
rect 293 2 356 9
rect 293 -63 315 2
rect 469 -2 490 64
rect 413 -10 490 -2
rect 413 -27 441 -10
rect 459 -27 490 -10
rect 413 -49 490 -27
rect 469 -61 490 -49
rect -62 -122 -42 -106
rect 29 -124 49 -106
rect 210 -123 232 -109
rect 293 -122 315 -109
rect 469 -120 490 -107
<< polycont >>
rect -226 7 -209 24
rect -90 7 -73 24
rect 0 12 18 29
rect 185 6 203 23
rect 321 9 339 26
rect 441 -27 459 -10
<< locali >>
rect 248 176 544 177
rect -118 175 544 176
rect -224 174 544 175
rect -224 173 189 174
rect -224 172 -179 173
rect -224 153 -216 172
rect -199 154 -179 172
rect -162 154 -145 173
rect -128 172 -36 173
rect -128 154 -97 172
rect -199 153 -97 154
rect -80 154 -36 172
rect -19 172 189 173
rect -19 154 62 172
rect -80 153 62 154
rect 79 155 189 172
rect 206 155 289 174
rect 306 155 376 174
rect 393 173 495 174
rect 393 156 431 173
rect 449 156 495 173
rect 393 155 495 156
rect 512 155 544 174
rect 79 153 544 155
rect -224 149 544 153
rect -224 148 -116 149
rect -220 108 -202 148
rect -236 98 -200 108
rect -236 70 -229 98
rect -209 70 -200 98
rect -236 60 -200 70
rect -179 100 -143 108
rect -93 104 -70 149
rect 62 104 81 149
rect 248 148 544 149
rect 153 107 210 108
rect 247 107 282 109
rect 322 107 360 108
rect 432 107 453 148
rect -179 72 -172 100
rect -152 72 -143 100
rect -179 60 -143 72
rect -105 97 -63 104
rect -105 69 -92 97
rect -72 69 -63 97
rect -105 61 -63 69
rect -30 98 6 103
rect -30 70 -22 98
rect -2 95 6 98
rect 1 78 6 95
rect -2 70 6 78
rect -30 62 6 70
rect 51 95 95 104
rect 51 67 60 95
rect 80 67 95 95
rect 51 61 95 67
rect 153 100 366 107
rect 153 97 253 100
rect 153 78 174 97
rect 198 78 253 97
rect 153 72 253 78
rect 273 95 366 100
rect 273 75 332 95
rect 350 76 366 95
rect 349 75 366 76
rect 273 72 366 75
rect 153 65 366 72
rect 426 96 463 107
rect 426 77 435 96
rect 452 77 463 96
rect 153 64 210 65
rect 247 64 282 65
rect -168 32 -150 60
rect -252 24 -201 30
rect -252 7 -226 24
rect -209 7 -201 24
rect -252 0 -201 7
rect -168 24 -63 32
rect -168 7 -90 24
rect -73 7 -63 24
rect -168 2 -63 7
rect -12 29 29 34
rect -12 12 0 29
rect 18 12 29 29
rect -12 3 29 12
rect 169 23 212 30
rect 169 6 185 23
rect 203 6 212 23
rect -168 -21 -150 2
rect 169 0 212 6
rect -92 -21 -66 -15
rect -238 -30 -200 -21
rect -238 -58 -231 -30
rect -211 -58 -200 -30
rect -238 -69 -200 -58
rect -179 -30 -143 -21
rect -179 -58 -172 -30
rect -152 -58 -143 -30
rect -179 -69 -143 -58
rect -92 -38 -86 -21
rect -69 -38 -66 -21
rect -92 -59 -66 -38
rect 249 -20 282 64
rect 322 63 360 65
rect 426 63 463 77
rect 498 96 535 108
rect 498 77 506 96
rect 523 77 535 96
rect 498 64 535 77
rect 310 26 356 33
rect 310 9 321 26
rect 339 9 356 26
rect 310 2 356 9
rect 506 5 530 64
rect 395 -10 475 -2
rect 249 -37 256 -20
rect 274 -37 282 -20
rect 249 -43 282 -37
rect 322 -18 355 -15
rect 395 -18 441 -10
rect 322 -20 441 -18
rect 322 -37 326 -20
rect 344 -27 441 -20
rect 459 -27 475 -10
rect 344 -37 475 -27
rect 322 -41 475 -37
rect 506 -24 579 5
rect -97 -69 -65 -59
rect -237 -145 -206 -69
rect -97 -97 -92 -69
rect -72 -97 -65 -69
rect -97 -105 -65 -97
rect 57 -73 89 -60
rect 57 -101 63 -73
rect 83 -101 89 -73
rect 57 -145 89 -101
rect 170 -72 202 -64
rect 322 -65 355 -41
rect 506 -61 530 -24
rect 170 -100 175 -72
rect 195 -100 202 -72
rect 170 -145 202 -100
rect 321 -78 355 -65
rect 321 -97 327 -78
rect 344 -97 355 -78
rect 321 -109 355 -97
rect 423 -70 459 -62
rect 423 -89 431 -70
rect 448 -89 459 -70
rect 423 -108 459 -89
rect 495 -75 531 -61
rect 495 -94 504 -75
rect 521 -94 531 -75
rect 495 -107 531 -94
rect 429 -143 452 -108
rect 252 -145 552 -143
rect -241 -149 552 -145
rect -241 -150 176 -149
rect -241 -153 60 -150
rect -241 -154 -180 -153
rect -241 -171 -233 -154
rect -216 -171 -180 -154
rect -241 -172 -180 -171
rect -163 -154 -14 -153
rect -163 -172 -102 -154
rect -241 -173 -102 -172
rect -85 -172 -14 -154
rect 3 -167 60 -153
rect 77 -166 176 -150
rect 193 -150 508 -149
rect 193 -166 240 -150
rect 77 -167 240 -166
rect 3 -169 240 -167
rect 257 -151 508 -150
rect 257 -152 432 -151
rect 257 -154 385 -152
rect 257 -169 327 -154
rect 3 -172 327 -169
rect -85 -173 327 -172
rect 344 -171 385 -154
rect 402 -168 432 -152
rect 449 -168 508 -151
rect 525 -168 552 -149
rect 402 -171 552 -168
rect 344 -173 552 -171
rect -241 -177 552 -173
rect 252 -178 552 -177
<< viali >>
rect -216 153 -199 172
rect -97 153 -80 172
rect 62 153 79 172
rect 431 156 449 173
rect -16 78 -2 95
rect -2 78 1 95
rect 174 78 181 97
rect 181 78 192 97
rect 332 94 350 95
rect 332 76 349 94
rect 349 76 350 94
rect -86 -38 -69 -21
rect 256 -37 274 -20
rect 326 -37 344 -20
rect -233 -171 -216 -154
rect 60 -167 77 -150
rect 176 -166 193 -149
rect 432 -168 449 -151
<< metal1 >>
rect 248 176 544 177
rect -118 175 544 176
rect -224 173 544 175
rect -224 172 431 173
rect -224 153 -216 172
rect -199 153 -97 172
rect -80 153 62 172
rect 79 156 431 172
rect 449 156 544 173
rect 79 153 544 156
rect -224 149 544 153
rect -224 148 -116 149
rect 248 148 544 149
rect 153 101 197 102
rect 153 99 364 101
rect -22 97 364 99
rect -22 95 174 97
rect -22 78 -16 95
rect 1 78 174 95
rect 192 95 364 97
rect 192 78 332 95
rect -22 76 332 78
rect 350 76 364 95
rect -22 75 212 76
rect 317 72 363 76
rect -92 -20 352 -16
rect -92 -21 256 -20
rect -92 -38 -86 -21
rect -69 -37 256 -21
rect 274 -37 326 -20
rect 344 -37 352 -20
rect -69 -38 352 -37
rect -92 -43 352 -38
rect 252 -145 552 -143
rect -241 -149 552 -145
rect -241 -150 176 -149
rect -241 -154 60 -150
rect -241 -171 -233 -154
rect -216 -167 60 -154
rect 77 -166 176 -150
rect 193 -151 552 -149
rect 193 -166 432 -151
rect 77 -167 432 -166
rect -216 -168 432 -167
rect 449 -168 552 -151
rect -216 -171 552 -168
rect -241 -177 552 -171
rect 252 -178 552 -177
<< labels >>
flabel locali -247 15 -247 15 0 FreeSans 80 0 0 0 s
port 2 nsew
flabel metal1 117 165 117 165 0 FreeSans 80 0 0 0 vdd
port 0 nsew
flabel polycont s 7 21 7 21 0 FreeSans 80 0 0 0 i0
port 4 nsew
flabel polycont s 178 20 178 20 0 FreeSans 80 0 0 0 i1
port 5 nsew
flabel polycont s 347 14 350 18 0 FreeSans 80 0 0 0 s
port 1 nsew
flabel locali s 541 -9 541 -9 0 FreeSans 80 0 0 0 y
port 7 nsew
flabel psubdiff s 112 -158 112 -158 0 FreeSans 80 0 0 0 gnd
port 9 nsew
<< end >>
