magic
tech scmos
timestamp 1735480075
<< nwell >>
rect -22 13 9 42
<< polysilicon >>
rect -10 25 -7 29
rect -10 -10 -7 17
rect -10 -20 -7 -15
<< ndiffusion >>
rect -12 -14 -10 -10
rect -17 -15 -10 -14
rect -7 -14 -4 -10
rect 1 -14 5 -10
rect -7 -15 5 -14
<< pdiffusion >>
rect -15 21 -10 25
rect -20 17 -10 21
rect -7 22 5 25
rect -7 18 -4 22
rect 1 18 5 22
rect -7 17 5 18
<< metal1 >>
rect -21 36 -17 41
rect -12 36 0 41
rect -20 25 -15 36
rect -4 5 1 18
rect -24 0 -17 4
rect -4 1 8 5
rect -4 -10 1 1
rect -17 -22 -12 -14
rect -18 -27 -15 -22
rect -10 -27 -3 -22
rect 2 -27 4 -22
<< ntransistor >>
rect -10 -15 -7 -10
<< ptransistor >>
rect -10 17 -7 25
<< polycontact >>
rect -17 0 -10 4
<< ndcontact >>
rect -17 -14 -12 -10
rect -4 -14 1 -10
<< pdcontact >>
rect -20 21 -15 25
rect -4 18 1 22
<< psubstratepcontact >>
rect -15 -27 -10 -22
rect -3 -27 2 -22
<< nsubstratencontact >>
rect -17 36 -12 41
rect 0 36 5 41
<< labels >>
rlabel metal1 -7 -24 -7 -24 1 gnd
rlabel metal1 8 3 8 3 7 out
rlabel metal1 -3 40 -3 40 5 vdd
rlabel metal1 -22 2 -22 2 3 in
<< end >>
