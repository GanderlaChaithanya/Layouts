* SPICE3 file created from inverter_design.ext - technology: scmos
.model pfet pmos level=49 version=3.3.0
.model nfet nmos level=49 version=3.3.0

.option scale=1u

M1000 out in vdd vdd pfet w=8 l=3
+  ad=96p pd=40u as=80p ps=36u
M1001 out in gnd Gnd nfet w=5 l=3
+  ad=60p pd=34u as=35p ps=24u
C0 gnd 0 4.47f **FLOATING
C1 out 0 6.72f **FLOATING
C2 in 0 14f **FLOATING

v1 vdd gnd 5
v1 in gnd pulse(0 5  0 1n 1n 10n 20n)

.tran 1n 100n
.control
run
plot V(in) V(out)

.endc
.end

