magic
tech sky130A
timestamp 1736604901
<< nwell >>
rect -159 -30 162 172
<< nmos >>
rect -79 -236 -40 -181
rect 42 -236 73 -181
<< pmos >>
rect -79 23 -40 77
rect 42 23 73 77
<< ndiff >>
rect -123 -195 -79 -181
rect -123 -221 -112 -195
rect -93 -221 -79 -195
rect -123 -236 -79 -221
rect -40 -236 42 -181
rect 73 -193 121 -181
rect 73 -219 84 -193
rect 103 -219 121 -193
rect 73 -236 121 -219
<< pdiff >>
rect -129 62 -79 77
rect -129 35 -117 62
rect -97 35 -79 62
rect -129 23 -79 35
rect -40 63 42 77
rect -40 36 -16 63
rect 4 36 42 63
rect -40 23 42 36
rect 73 63 124 77
rect 73 31 86 63
rect 111 31 124 63
rect 73 23 124 31
<< ndiffc >>
rect -112 -221 -93 -195
rect 84 -219 103 -193
<< pdiffc >>
rect -117 35 -97 62
rect -16 36 4 63
rect 86 31 111 63
<< psubdiff >>
rect -130 -300 155 -295
rect -130 -301 14 -300
rect -130 -327 -105 -301
rect -80 -326 14 -301
rect 39 -326 155 -300
rect -80 -327 155 -326
rect -130 -332 155 -327
<< nsubdiff >>
rect -141 150 130 154
rect -141 149 15 150
rect -141 122 -53 149
rect -30 123 15 149
rect 38 123 130 150
rect -30 122 130 123
rect -141 117 130 122
<< psubdiffcont >>
rect -105 -327 -80 -301
rect 14 -326 39 -300
<< nsubdiffcont >>
rect -53 122 -30 149
rect 15 123 38 150
<< poly >>
rect -79 77 -40 99
rect 42 77 73 97
rect -79 -54 -40 23
rect -138 -61 -40 -54
rect -138 -83 -119 -61
rect -96 -83 -40 -61
rect -138 -89 -40 -83
rect -79 -181 -40 -89
rect 42 -39 73 23
rect 42 -47 110 -39
rect 42 -69 79 -47
rect 102 -69 110 -47
rect 42 -78 110 -69
rect 42 -181 73 -78
rect -79 -270 -40 -236
rect 42 -275 73 -236
<< polycont >>
rect -119 -83 -96 -61
rect 79 -69 102 -47
<< locali >>
rect -132 154 126 155
rect -141 150 126 154
rect -141 149 15 150
rect -141 148 -53 149
rect -141 121 -119 148
rect -96 122 -53 148
rect -30 123 15 149
rect 38 149 126 150
rect 38 123 87 149
rect -30 122 87 123
rect 110 122 126 149
rect -96 121 126 122
rect -141 117 126 121
rect -124 62 -91 117
rect -124 35 -117 62
rect -97 35 -91 62
rect -124 27 -91 35
rect -21 63 9 71
rect -21 36 -16 63
rect 4 36 9 63
rect -161 -61 -79 -54
rect -161 -83 -119 -61
rect -96 -83 -79 -61
rect -161 -90 -79 -83
rect -117 -119 -85 -115
rect -117 -143 -112 -119
rect -91 -143 -85 -119
rect -117 -195 -85 -143
rect -21 -118 9 36
rect 79 70 121 117
rect 79 63 120 70
rect 79 31 86 63
rect 111 31 120 63
rect 79 23 120 31
rect 73 -47 144 -39
rect 73 -69 79 -47
rect 102 -69 144 -47
rect 73 -78 144 -69
rect -21 -142 -17 -118
rect 4 -142 9 -118
rect -21 -145 9 -142
rect -117 -221 -112 -195
rect -93 -221 -85 -195
rect -117 -229 -85 -221
rect 76 -193 111 -186
rect 76 -219 84 -193
rect 103 -219 111 -193
rect 76 -295 111 -219
rect -130 -300 155 -295
rect -130 -301 14 -300
rect -130 -327 -105 -301
rect -80 -326 14 -301
rect 39 -301 155 -300
rect 39 -326 81 -301
rect -80 -327 81 -326
rect 106 -327 155 -301
rect -130 -332 155 -327
rect 76 -333 111 -332
<< viali >>
rect -119 121 -96 148
rect 87 122 110 149
rect -112 -143 -91 -119
rect -17 -142 4 -118
rect 81 -327 106 -301
<< metal1 >>
rect -140 149 126 154
rect -140 148 87 149
rect -140 121 -119 148
rect -96 122 87 148
rect 110 122 126 149
rect -96 121 126 122
rect -140 117 126 121
rect -151 -118 119 -115
rect -151 -119 -17 -118
rect -151 -143 -112 -119
rect -91 -142 -17 -119
rect 4 -142 119 -118
rect -91 -143 119 -142
rect -151 -146 119 -143
rect -126 -301 153 -295
rect -126 -327 81 -301
rect 106 -327 153 -301
rect -126 -333 153 -327
<< labels >>
flabel metal1 -11 135 -11 135 0 FreeSans 80 0 0 0 vdd
flabel metal1 -33 -320 -33 -320 0 FreeSans 80 0 0 0 gnd
flabel locali -149 -74 -149 -74 0 FreeSans 160 0 0 0 A
flabel locali 122 -62 122 -62 0 FreeSans 160 0 0 0 B
flabel metal1 93 -129 93 -129 0 FreeSans 160 0 0 0 OUT
<< end >>
